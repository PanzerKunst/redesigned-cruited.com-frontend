# Global

signIn=Sign in

product.name.CV_REVIEW=CV [Resume]
product.name.COVER_LETTER_REVIEW=Cover Letter
product.name.LINKEDIN_PROFILE_REVIEW=Linkedin Profile

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive

reduction.name.2_PRODUCTS_SAME_ORDER=2-item
reduction.name.3_PRODUCTS_SAME_ORDER=3-item


# Order Step Product Selection page

orderStepProductSelection.title=Product Selection
orderStepProductSelection.subtitle=How can we help you?
orderStepProductSelection.nextStepBtn.text=Proceed to next step

orderStepProductSelection.productsSection.title=Products
orderStepProductSelection.productsSection.offerTwoProductsSameOrder.text=Save <strong>{reductionPrice}</strong> off your order when you select 2 items!
orderStepProductSelection.productsSection.offerThreeProductsSameOrder.text=Save <strong>{reductionPrice}</strong> off your order when you select all 3 items!
orderStepProductSelection.productsSection.productName.CV_REVIEW=Review my CV
orderStepProductSelection.productsSection.productName.COVER_LETTER_REVIEW=Review my Cover Letter
orderStepProductSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Review my Linkedin Profile

orderStepProductSelection.editionsSection.title=Product Edition
orderStepProductSelection.editionsSection.subtitle=Please choose which edition best suits you

orderStepProductSelection.cartSection.title=Your Order
orderStepProductSelection.cartSection.productsHeader.products=Products
orderStepProductSelection.cartSection.productsHeader.defaultPrice=Price
orderStepProductSelection.cartSection.edition=Edition
orderStepProductSelection.cartSection.coupon.label=Have a valid Promotion code or a Gift Card from one of our partners?
orderStepProductSelection.cartSection.coupon.field.placeholder=Coupon Code
orderStepProductSelection.cartSection.coupon.addBtn.text=Apply coupon
orderStepProductSelection.cartSection.coupon.addBtn.loadingText=Applying coupon...
orderStepProductSelection.cartSection.coupon.notFoundError=Coupon not found or expired
orderStepProductSelection.cartSection.subTotal=Sub-total
orderStepProductSelection.cartSection.total=Total You Pay


# Order Step AssessmentInfo page

orderStepAssessmentInfo.title=Assessment details
orderStepAssessmentInfo.subtitle=Tell us a bit about you
orderStepAssessmentInfo.nextStepBtn.text=Proceed to next step

orderStepAssessmentInfo.form.field.browseBtn.text=Browse...
orderStepAssessmentInfo.form.field.linkedinProfile.label=Your Linkedin profile
orderStepAssessmentInfo.form.field.linkedinProfile.signInBtn.text=Sign in with Linkedin
orderStepAssessmentInfo.form.field.linkedinProfile.check.step1.text=Öppna nu <a href="https://www.linkedin.com/profile/public-profile-settings?trk=prof-edit-edit-public_profile" target="blank">dina profilinställningar</a> och se till att alla kryssrutor till höger är ifyllda. De delar du inte kryssar för kommer vi inte att kunna granska.
orderStepAssessmentInfo.form.field.linkedinProfile.check.step2.text=Ta en titt på <a href="https://www.linkedin.com/profile/preview?vpa=pub" target="blank">din publika profilsida</a> och se till att all information är synlig. Det du ser här är det vi kommer att bedöma.
orderStepAssessmentInfo.form.field.linkedinProfile.check.checkbox.label=Klart! Min profil är redo för granskning
orderStepAssessmentInfo.form.field.linkedinProfile.validation.notSignedIn=We cannot assess your Linkedin profile unless you sign in
orderStepAssessmentInfo.form.field.cvFile.label=Your CV
orderStepAssessmentInfo.form.field.cvFile.placeHolder=PDF, Word, ...
orderStepAssessmentInfo.form.field.coverLetterFile.label=Your cover letter
orderStepAssessmentInfo.form.field.coverLetterFile.placeHolder=PDF, Word, ...
orderStepAssessmentInfo.form.field.employerSought.label=Employer sought
orderStepAssessmentInfo.form.field.positionSought.label=Position sought
orderStepAssessmentInfo.form.field.jobAdUrl.label=URL of the job ad
orderStepAssessmentInfo.form.tos.text=I have read and accept the <a>Terms of Service</a>
