# Global

defaultAssessmentTitle=

product.name.CV_REVIEW=Granskning av CV
product.name.COVER_LETTER_REVIEW=Granskning av personligt brev
product.name.LINKEDIN_PROFILE_REVIEW=Granskning av LinkedIn

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive
edition.name.short.PRO=Professional
edition.name.short.YOUNG_PRO=Young Pro
edition.name.short.EXEC=Executive

reduction.name.2_PRODUCTS_SAME_ORDER=2 dokument
reduction.name.3_PRODUCTS_SAME_ORDER=3 dokument

order.status.label=Status
order.status.notPaid.text=Betalning saknas
order.status.paid.text=Avvaktar granskning
order.status.inProgress.text=Granskning pågår
order.status.completed.text=Granskning genomförd

order.creationDate.label=Skapad

category.CV_REVIEW.12.title=Redovisa resultat och skapa trovärdighet
category.CV_REVIEW.12.shortDesc=En cv handlar i stor utsträckning om att bekräfta sin kompetens. Det är därför mycket viktigt att redovisa de resultat man uppnått.
category.CV_REVIEW.13.title=Översiktligt och korrekt
category.CV_REVIEW.13.shortDesc=Din cv ska ge arbetsgivaren en snabb översikt över dina erfarenheter och meriter. Den ska vara korrekt skriven, kort och koncis. Det finns även ett antal faktorer i språk och upplägget som påverkar hur du uppfattas som person.
category.CV_REVIEW.14.title=Rikta och var relevant
category.CV_REVIEW.14.shortDesc=I en effektiv cv är varje del relevant för det aktuella jobbet och den aktuella arbetsgivaren. Det kräver att cvn har en tydlig röd linje och att alla delar pekar i samma riktning.
category.COVER_LETTER_REVIEW.7.title=Framhäv potential
category.COVER_LETTER_REVIEW.7.shortDesc=Fokusera mer på din potential och vad du kan åstadkomma i framtiden, än på historia och vad du gjort tidigare.
category.COVER_LETTER_REVIEW.8.title=Fokusera på arbetsgivaren
category.COVER_LETTER_REVIEW.8.shortDesc=Förklara varför du valt just den här arbetsgivaren och tjänsten.
category.COVER_LETTER_REVIEW.10.title=Redovisa resultat och skapa trovärdighet
category.COVER_LETTER_REVIEW.10.shortDesc=Visa på ett trovärdigt sätt att du har kunskapen och förmågan att åstadkomma resultat för arbetsgivaren.
category.COVER_LETTER_REVIEW.11.title=Aktivt, kort och korrekt
category.COVER_LETTER_REVIEW.11.shortDesc=En dåligt skriven ansökan placerar dig som sökande ofta direkt längst ner i högen.
category.LINKEDIN_PROFILE_REVIEW.16.title=Rikta och var relevant
category.LINKEDIN_PROFILE_REVIEW.16.shortDesc=Nyckeln till framgång bland miljontals profiler på LinkedIn är att vara relevant. Du behöver visa en röd linje, få fram en bild av vart du är på väg och vad du söker. I vår granskning tittar vi på flera faktorer som rör relevans och riktning.
category.LINKEDIN_PROFILE_REVIEW.17.title=Skapa effekt och bygg räckvidd
category.LINKEDIN_PROFILE_REVIEW.17.shortDesc=Att finnas på LinkedIn är grundläggande när man söker jobb. Men för att nå framgång med LinkedIn behöver man synas och underlätta kontaktskapande. Den här kategorin handlar om hur du lyckas skapa effekt och nå ut med din profil.
category.LINKEDIN_PROFILE_REVIEW.18.title=Översiktligt och korrekt
category.LINKEDIN_PROFILE_REVIEW.18.shortDesc=Din LinkedIn-profil ska vara korrekt skriven och lätt att ta till sig. För att bli hittad av rekryterare och andra som vill nå dig, är det också viktigt att profilen är komplett och att du fyllt i rätt uppgifter på rätt plats.
category.LINKEDIN_PROFILE_REVIEW.20.title=Redovisa resultat och skapa trovärdighet
category.LINKEDIN_PROFILE_REVIEW.20.shortDesc=LinkedIn är världens största cv-bank och att berätta om sina erfarenheter och utbildningar är grundläggande. För att få kontakter och skapa möjligheter till jobb behöver du ge trovärdig bild av din bakgrund.

reportSummary.CV_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du har en bra bit kvar innan vi kan rekommendera dig att skicka in denna jobbansökan. Läs gärna våra rekommendationer nedan för att göra en mer genomarbetad version av din CV. Du har möjligheten att göra en stor förbättring ganska lätt om du följer dem!
reportSummary.CV_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du borde göra ett nytt försök, för du har en bit kvar innan du har skrivit en jobbansökan som du med stolthet kan skicka in till din potentiella arbetsgivare. Följ gärna våra rekommendationer nedan för att få din ansökan att hålla den klass vi tror att du vill att den ska hålla!
reportSummary.CV_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du har gjort en bra insats, det är helt okej, men du borde jobba vidare med din jobbansökan. Följ gärna våra rekommendationer nedan så kan din ansökan bli exemplariskt bra!
reportSummary.CV_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du kan vara mycket nöjd med din insats! Överväg gärna att följa våra råd till förbättringar nedan - du är inte många steg ifrån att ha gjort en utmärkt jobbansökan!
reportSummary.CV_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Mycket bra jobbat! Ditt ansökningsbrev är riktigt riktigt bra! Det skadar förstås aldrig att ändå ta en titt på råden nedan för att se om det är något du kan förbättra ytterligare. Men var stolt över din insats!
reportSummary.COVER_LETTER_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du har en bra bit kvar innan vi kan rekommendera dig att skicka in denna jobbansökan. Läs gärna våra rekommendationer nedan för att göra en mer genomarbetad version av ditt personliga brev. Du har möjligheten att göra en stor förbättring ganska lätt om du följer dem!
reportSummary.COVER_LETTER_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du borde göra ett nytt försök, för du har en bit kvar innan du har skrivit en jobbansökan som du med stolthet kan skicka in till din potentiella arbetsgivare. Följ gärna våra rekommendationer nedan för att få din ansökan att hålla den klass vi tror att du vill att den ska hålla!
reportSummary.COVER_LETTER_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du har gjort en bra insats, det är helt okej, men du borde jobba vidare med din jobbansökan. Följ gärna våra rekommendationer nedan så kan din ansökan bli exemplariskt bra!
reportSummary.COVER_LETTER_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du kan vara mycket nöjd med din insats! Överväg gärna att följa våra råd till förbättringar nedan - du är inte många steg ifrån att ha gjort en utmärkt jobbansökan!
reportSummary.COVER_LETTER_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Mycket bra jobbat! Ditt ansökningsbrev är riktigt riktigt bra! Det skadar förstås aldrig att ändå ta en titt på råden nedan för att se om det är något du kan förbättra ytterligare. Men var stolt över din insats!
reportSummary.LINKEDIN_PROFILE_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din Linkedin-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av Linkedin-profil är <strong>{averageScore}</strong>.<br /><br />Du har en bra bit kvar innan du har en profil som kommer att locka rekryterare och potentiella arbetsgivare. Läs gärna våra rekommendationer nedan för att göra en mer genomarbetad version av din Linkedin-profil. Du har möjligheten att göra en stor förbättring ganska lätt om du följer dem!
reportSummary.LINKEDIN_PROFILE_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din Linkedin-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av Linkedin-profil är <strong>{averageScore}</strong>.<br /><br />Du borde göra ett nytt försök, för du har en bit kvar innan du har en profil som sticker ut hos en rekryterare eller potentiell arbetsgivare. Följ gärna våra rekommendationer nedan för att få din profil att hålla den klass vi tror att du vill att den ska hålla!
reportSummary.LINKEDIN_PROFILE_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din Linkedin-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av Linkedin-profil är <strong>{averageScore}</strong>.<br /><br />Du har gjort en bra insats, det är helt okej, men du borde jobba vidare med din profil. Följ gärna våra rekommendationer nedan så kan din profil bli exemplariskt bra!
reportSummary.LINKEDIN_PROFILE_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din Linkedin-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av Linkedin-profil är <strong>{averageScore}</strong>.<br /><br />Du kan vara mycket nöjd med din insats! Överväg gärna att följa våra råd till förbättringar nedan - du är inte många steg ifrån att ha gjort en utmärkt profil!
reportSummary.LINKEDIN_PROFILE_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din Linkedin-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av Linkedin-profil är <strong>{averageScore}</strong>.<br /><br />Mycket bra jobbat! Din profil är riktigt riktigt bra! Det skadar förstås aldrig att ändå ta en titt på råden nedan för att se om det är något du kan förbättra ytterligare. Men var stolt över din insats!


# Header menu

menu.signIn=Logga in
menu.signOut=Logga ut
menu.myAccount=Mitt konto


# Sign In page

signIn.title=Logga in
signIn.methodSeparatorText=eller...
signIn.validation.incorrectEmail=Den här e-postadressen ser inte korrekt ut
signIn.validation.invalidCredentials=Vi har inget konto med den här adressen
signIn.validation.linkedinAccountUnregistered=Du har inget konto kopplat till den här Linkedin . Registrera dig Registration is done during <a href="/order">your first order</a>.

signIn.form.linkedIn.btn.text=
signIn.form.email.emailAddress.label=
signIn.form.email.emailAddress.placeholder=
signIn.form.email.password.label=
signin.form.email.submitBtn.text=
signIn.form.forgottenPasswordLink.text=


# My Account page

myAccount.title=
myAccount.validation.passwordTooShort=
myAccount.saveSuccessful.text=

myAccount.form.emailAddress.label=
myAccount.form.firstName.label=
myAccount.form.password.label=
myAccount.form.password.placeholder=
myAccount.form.submitBtn.text=


# Reset password pages

resetPassword.title=
resetPassword.validation.incorrectEmail=
resetPassword.validation.noAccountFoundForThisEmailAddress=
resetPassword.emailSent.text=

resetPassword.form.emailAddress.label=
resetPassword.form.emailAddress.placeholder=
resetPassword.form.submitBtn.text=

resetPassword.new.saveSuccessful.text=
resetPassword.new.validation.passwordTooShort=
resetPassword.new.form.password.label=
resetPassword.new.form.password.placeholder=
resetPassword.new.form.submitBtn.text=


# Dashboard page

dashboard.title=
dashboard.subtitle=
dashboard.completePaymentLink.text=
dashboard.newAssessmentBtn.text=
dashboard.viewReportBtn.text=
dashboard.editOrder.text=


# Report page

report.title=
report.unorderedAssessment.text=
report.unorderedAssessment.orderBtn.text=

report.summary.title=
report.summary.documentLink.text=
report.summary.score.label=
report.summary.score.bar.label.weak=
report.summary.score.bar.label.good=
report.summary.score.bar.label.excellent=
report.summary.understandYourScore.title=
report.summary.understandYourScore.cScoreExplanation.text=
report.summary.understandYourScore.weak.text=
report.summary.understandYourScore.good.text=
report.summary.understandYourScore.excellent.text=

report.analysis.title=


# Order Step Product Selection page

order.productSelection.title=
order.productSelection.subtitle=
order.productSelection.submitBtn.text=
order.productSelection.validation.emptyCart=

order.productSelection.productsSection.title=
order.productSelection.productsSection.offerTwoProductsSameOrder.text=
order.productSelection.productsSection.offerThreeProductsSameOrder.text=
order.productSelection.productsSection.allOffersActivated.text=
order.productSelection.productsSection.productName.CV_REVIEW=
order.productSelection.productsSection.productName.COVER_LETTER_REVIEW=
order.productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=

order.productSelection.editionsSection.title=
order.productSelection.editionsSection.subtitle=
order.productSelection.editionsSection.editionDescription.text.PRO=
order.productSelection.editionsSection.editionDescription.text.YOUNG_PRO=
order.productSelection.editionsSection.editionDescription.text.EXEC=

order.productSelection.cartSection.title=
order.productSelection.cartSection.productsHeader.products=
order.productSelection.cartSection.productsHeader.defaultPrice=
order.productSelection.cartSection.coupon.label=
order.productSelection.cartSection.coupon.placeholder=
order.productSelection.cartSection.coupon.addBtn.text=
order.productSelection.cartSection.coupon.addBtn.loadingText=
order.productSelection.cartSection.coupon.notFoundError=
order.productSelection.cartSection.coupon.hasReachedMaxUsesError=
order.productSelection.cartSection.subTotal=
order.productSelection.cartSection.total=


# Order Step Assessment Info page

order.assessmentInfo.title=
order.assessmentInfo.subtitle=
order.assessmentInfo.documentsSection.title=
order.assessmentInfo.documentsSection.subtitle=
order.assessmentInfo.jobYouSearchSection.title=
order.assessmentInfo.jobYouSearchSection.subtitle=
order.assessmentInfo.submitBtn.text=
order.assessmentInfo.validation.notSignedIn=
order.assessmentInfo.validation.jobAdUrlIncorrect=
order.assessmentInfo.validation.customerCommentTooLong=

order.assessmentInfo.form.browseBtn.text=
order.assessmentInfo.form.linkedinProfile.label=
order.assessmentInfo.form.linkedinProfile.signInBtn.text=
order.assessmentInfo.form.linkedinProfile.check.step1.text=
order.assessmentInfo.form.linkedinProfile.check.step2.text=
order.assessmentInfo.form.linkedinProfile.check.checkbox.label=
order.assessmentInfo.form.cvFile.label=
order.assessmentInfo.form.cvFile.placeHolder=
order.assessmentInfo.form.coverLetterFile.label=
order.assessmentInfo.form.coverLetterFile.placeHolder=
order.assessmentInfo.form.employerSought.label=
order.assessmentInfo.form.positionSought.label=
order.assessmentInfo.form.jobAdUrl.label=
order.assessmentInfo.form.customerComment.label=
order.assessmentInfo.form.customerComment.description=
order.assessmentInfo.form.tos.text=


# Order Step Account Creation page

order.accountCreation.title=
order.accountCreation.subtitle=
order.accountCreation.submitBtn.text=
order.accountCreation.submitBtn.withEmailPrefix=
order.accountCreation.validation.emailAlreadyRegistered=
order.accountCreation.validation.linkedinAccountIdAlreadyRegistered=

order.accountCreation.registerWithLinkedin.switchLink.text=
order.accountCreation.registerWithLinkedin.btn.text=
order.accountCreation.registerWithLinkedin.email.label=
order.accountCreation.registerWithLinkedin.validation.incorrectEmail=

order.accountCreation.registerWithEmail.switchLink.text=
order.accountCreation.registerWithEmail.firstName.label=
order.accountCreation.registerWithEmail.firstName.placeholder=
order.accountCreation.registerWithEmail.emailAddress.label=
order.accountCreation.registerWithEmail.emailAddress.placeholder=
order.accountCreation.registerWithEmail.password.label=
order.accountCreation.registerWithEmail.password.placeholder=
order.accountCreation.registerWithEmail.validation.incorrectEmail=
order.accountCreation.registerWithEmail.validation.passwordTooShort=


# Order Step Payment page

order.payment.title=
order.payment.subtitle=
order.payment.submitBtn.text=
order.payment.validation.invalidCardNumber=
order.payment.validation.invalidExpirationDate=
order.payment.success.text=

order.payment.form.cardNumber.label=
order.payment.form.cardNumber.placeholder=
order.payment.form.expires.month.label=
order.payment.form.cvc.label=
order.payment.form.cvc.placeholder=
order.payment.form.cardholderName.label=


# Edit Order page

order.edit.saveBtn.text=


# Emails

email.resetPassword.subject=
email.unpaidOrderReminder.subject=
email.twoDaysAfterAssessmentDelivered.subject=
email.orderComplete.free.subject=
email.orderComplete.paid.subject=
email.orderComplete.paid.orderedProductsSeparator=
