# Global

defaultAssessmentTitle=Bedömning

product.name.CV_REVIEW=Granskning av CV
product.name.COVER_LETTER_REVIEW=Granskning av personligt brev
product.name.LINKEDIN_PROFILE_REVIEW=Granskning av LinkedIn

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive
edition.name.short.PRO=Professional
edition.name.short.YOUNG_PRO=Young Pro
edition.name.short.EXEC=Executive

reduction.name.2_PRODUCTS_SAME_ORDER=2 dokument
reduction.name.3_PRODUCTS_SAME_ORDER=3 dokument

order.status.label=Status
order.status.notPaid.text=Betalning saknas
order.status.paid.text=Avvaktar granskning
order.status.inProgress.text=Granskning pågår
order.status.completed.text=Granskning genomförd

order.creationDate.label=Skapad

category.CV_REVIEW.12.title=Redovisa resultat och skapa trovärdighet
category.CV_REVIEW.12.shortDesc=En cv handlar i stor utsträckning om att bekräfta sin kompetens. Det är därför mycket viktigt att redovisa de resultat man uppnått.
category.CV_REVIEW.13.title=Översiktligt och korrekt
category.CV_REVIEW.13.shortDesc=Din cv ska ge arbetsgivaren en snabb översikt över dina erfarenheter och meriter. Den ska vara korrekt skriven, kort och koncis. Det finns även ett antal faktorer i språk och upplägget som påverkar hur du uppfattas som person.
category.CV_REVIEW.14.title=Rikta och var relevant
category.CV_REVIEW.14.shortDesc=I en effektiv cv är varje del relevant för det aktuella jobbet och den aktuella arbetsgivaren. Det kräver att cvn har en tydlig röd linje och att alla delar pekar i samma riktning.
category.COVER_LETTER_REVIEW.7.title=Framhäv potential
category.COVER_LETTER_REVIEW.7.shortDesc=Fokusera mer på din potential och vad du kan åstadkomma i framtiden, än på historia och vad du gjort tidigare.
category.COVER_LETTER_REVIEW.8.title=Fokusera på arbetsgivaren
category.COVER_LETTER_REVIEW.8.shortDesc=Förklara varför du valt just den här arbetsgivaren och tjänsten.
category.COVER_LETTER_REVIEW.10.title=Redovisa resultat och skapa trovärdighet
category.COVER_LETTER_REVIEW.10.shortDesc=Visa på ett trovärdigt sätt att du har kunskapen och förmågan att åstadkomma resultat för arbetsgivaren.
category.COVER_LETTER_REVIEW.11.title=Aktivt, kort och korrekt
category.COVER_LETTER_REVIEW.11.shortDesc=En dåligt skriven ansökan placerar dig som sökande ofta direkt längst ner i högen.
category.LINKEDIN_PROFILE_REVIEW.16.title=Rikta och var relevant
category.LINKEDIN_PROFILE_REVIEW.16.shortDesc=Nyckeln till framgång bland miljontals profiler på LinkedIn är att vara relevant. Du behöver visa en röd linje, få fram en bild av vart du är på väg och vad du söker. I vår granskning tittar vi på flera faktorer som rör relevans och riktning.
category.LINKEDIN_PROFILE_REVIEW.17.title=Skapa effekt och bygg räckvidd
category.LINKEDIN_PROFILE_REVIEW.17.shortDesc=Att finnas på LinkedIn är grundläggande när man söker jobb. Men för att nå framgång med LinkedIn behöver man synas och underlätta kontaktskapande. Den här kategorin handlar om hur du lyckas skapa effekt och nå ut med din profil.
category.LINKEDIN_PROFILE_REVIEW.18.title=Översiktligt och korrekt
category.LINKEDIN_PROFILE_REVIEW.18.shortDesc=Din LinkedIn-profil ska vara korrekt skriven och lätt att ta till sig. För att bli hittad av rekryterare och andra som vill nå dig, är det också viktigt att profilen är komplett och att du fyllt i rätt uppgifter på rätt plats.
category.LINKEDIN_PROFILE_REVIEW.20.title=Redovisa resultat och skapa trovärdighet
category.LINKEDIN_PROFILE_REVIEW.20.shortDesc=LinkedIn är världens största cv-bank och att berätta om sina erfarenheter och utbildningar är grundläggande. För att få kontakter och skapa möjligheter till jobb behöver du ge trovärdig bild av din bakgrund.

reportSummary.CV_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du har en bra bit kvar innan vi kan rekommendera dig att skicka in denna jobbansökan. Läs gärna våra rekommendationer nedan för att göra en mer genomarbetad version av din CV. Du har möjligheten att göra en stor förbättring ganska lätt om du följer dem!
reportSummary.CV_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du borde göra ett nytt försök, för du har en bit kvar innan du har skrivit en jobbansökan som du med stolthet kan skicka in till din potentiella arbetsgivare. Följ gärna våra rekommendationer nedan för att få din ansökan att hålla den klass vi tror att du vill att den ska hålla!
reportSummary.CV_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du har gjort en bra insats, det är helt okej, men du borde jobba vidare med din jobbansökan. Följ gärna våra rekommendationer nedan så kan din ansökan bli exemplariskt bra!
reportSummary.CV_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Du kan vara mycket nöjd med din insats! Överväg gärna att följa våra råd till förbättringar nedan - du är inte många steg ifrån att ha gjort en utmärkt jobbansökan!
reportSummary.CV_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista CV granskningarna är <strong>{averageScore}</strong>.<br /><br />Mycket bra jobbat! Ditt ansökningsbrev är riktigt riktigt bra! Det skadar förstås aldrig att ändå ta en titt på råden nedan för att se om det är något du kan förbättra ytterligare. Men var stolt över din insats!
reportSummary.COVER_LETTER_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du har en bra bit kvar innan vi kan rekommendera dig att skicka in denna jobbansökan. Läs gärna våra rekommendationer nedan för att göra en mer genomarbetad version av ditt personliga brev. Du har möjligheten att göra en stor förbättring ganska lätt om du följer dem!
reportSummary.COVER_LETTER_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du borde göra ett nytt försök, för du har en bit kvar innan du har skrivit en jobbansökan som du med stolthet kan skicka in till din potentiella arbetsgivare. Följ gärna våra rekommendationer nedan för att få din ansökan att hålla den klass vi tror att du vill att den ska hålla!
reportSummary.COVER_LETTER_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du har gjort en bra insats, det är helt okej, men du borde jobba vidare med din jobbansökan. Följ gärna våra rekommendationer nedan så kan din ansökan bli exemplariskt bra!
reportSummary.COVER_LETTER_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Du kan vara mycket nöjd med din insats! Överväg gärna att följa våra råd till förbättringar nedan - du är inte många steg ifrån att ha gjort en utmärkt jobbansökan!
reportSummary.COVER_LETTER_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av personligt brev är <strong>{averageScore}</strong>.<br /><br />Mycket bra jobbat! Ditt ansökningsbrev är riktigt riktigt bra! Det skadar förstås aldrig att ändå ta en titt på råden nedan för att se om det är något du kan förbättra ytterligare. Men var stolt över din insats!
reportSummary.LINKEDIN_PROFILE_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.<br /><br />Du har en bra bit kvar innan du har en profil som kommer att locka rekryterare och potentiella arbetsgivare. Läs gärna våra rekommendationer nedan för att göra en mer genomarbetad version av din LinkedIn-profil. Du har möjligheten att göra en stor förbättring ganska lätt om du följer dem!
reportSummary.LINKEDIN_PROFILE_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.<br /><br />Du borde göra ett nytt försök, för du har en bit kvar innan du har en profil som sticker ut hos en rekryterare eller potentiell arbetsgivare. Följ gärna våra rekommendationer nedan för att få din profil att hålla den klass vi tror att du vill att den ska hålla!
reportSummary.LINKEDIN_PROFILE_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.<br /><br />Du har gjort en bra insats, det är helt okej, men du borde jobba vidare med din profil. Följ gärna våra rekommendationer nedan så kan din profil bli exemplariskt bra!
reportSummary.LINKEDIN_PROFILE_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.<br /><br />Du kan vara mycket nöjd med din insats! Överväg gärna att följa våra råd till förbättringar nedan - du är inte många steg ifrån att ha gjort en utmärkt profil!
reportSummary.LINKEDIN_PROFILE_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} sista granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.<br /><br />Mycket bra jobbat! Din profil är riktigt riktigt bra! Det skadar förstås aldrig att ändå ta en titt på råden nedan för att se om det är något du kan förbättra ytterligare. Men var stolt över din insats!


# Header menu

menu.signIn=Logga in
menu.signOut=Logga ut
menu.myAccount=Mitt konto


# Footer


# Sign In page

signIn.title=Logga in
signIn.methodSeparatorText=eller
signIn.validation.incorrectEmail=Den här e-postadressen ser inte korrekt ut
signIn.validation.invalidCredentials=Vi har inget konto med den här adressen
signIn.validation.linkedinAccountUnregistered=Vi kunde inte hitta ett konto hos oss kopplat till ditt på LinkedIn. Du kanske registrerade dig hos oss med din e-postadress? 

signIn.form.linkedIn.btn.text=Logga in med LinkedIn
signIn.form.email.emailAddress.label=E-postadress
signIn.form.email.emailAddress.placeholder=din@e-post.com
signIn.form.email.password.label=Lösenord
signin.form.email.submitBtn.text=Logga in
signIn.form.forgottenPasswordLink.text=Jag behöver ett nytt lösenord


# My Account page

myAccount.title=Mitt konto
myAccount.validation.passwordTooShort=Lösenordet behöver vara minst 5 tecken
myAccount.saveSuccessful.text=Ditt konto har uppdaterats

myAccount.form.emailAddress.label=E-postadress
myAccount.form.firstName.label=Förnamn
myAccount.form.password.label=Nytt lösenord (bara om du vill byta)
myAccount.form.password.placeholder=Minst 5 tecken
myAccount.form.submitBtn.text=Spara


# Reset password pages

resetPassword.title=Återställ ditt lösenord
resetPassword.validation.incorrectEmail=Den här e-postadressen ser inte korrekt ut
resetPassword.validation.noAccountFoundForThisEmailAddress=Vi har inget konto med den här adressen
resetPassword.emailSent.text=Vi har skickat ett mejl till dig med instruktioner om hur du återställer ditt lösenord

resetPassword.form.emailAddress.label=E-postadress
resetPassword.form.emailAddress.placeholder=din@e-post.com
resetPassword.form.submitBtn.text=Jag behöver ett nytt lösenord

resetPassword.new.saveSuccessful.text=Ditt nya lösenord är sparat. Nu kan du <a href="/login">logga in</a>.
resetPassword.new.validation.passwordTooShort=Lösenordet behöver vara minst 5 tecken
resetPassword.new.form.password.label=Nytt lösenord
resetPassword.new.form.password.placeholder=Minst 5 tecken
resetPassword.new.form.submitBtn.text=Spara


# Dashboard page

dashboard.title=Mina granskningar
dashboard.subtitle=Välkommen, {firstName}!
dashboard.completePaymentLink.text=Betala
dashboard.newAssessmentBtn.text=Skapa ny granskning
dashboard.viewReportBtn.text=Visa rapport
dashboard.editOrder.text=Den här granskningen har inte påbörjats och du kan fortfarande <a href="{url}">redigera din information</a> om du vill.


# Report page

report.title=Your Report
report.unorderedAssessment.text=You have not ordered this product. If you want to proceed, please place a new order.
report.unorderedAssessment.orderBtn.text=Order a new assessment
report.tabNameSmallScreen.CV_REVIEW=CV
report.tabNameSmallScreen.COVER_LETTER_REVIEW=Cover Letter
report.tabNameSmallScreen.LINKEDIN_PROFILE_REVIEW=LinkedIn

report.summary.title=Analysis of your document
report.summary.documentLink.text=Original doc
report.summary.score.label=Your C-Score
report.summary.score.bar.label.weak=Weak
report.summary.score.bar.label.good=Good
report.summary.score.bar.label.excellent=Excellent
report.summary.understandYourScore.title=Understand your score
report.summary.understandYourScore.cScoreExplanation.text=C-Score mäter hur effektiv din ansökan är på en skala från 0 till 100. <a href="https://www.cruited.com/var-metod" target="_blank">Läs mer</a>
report.summary.understandYourScore.weak.text=Mycket låg chans att komma på jobbintervju
report.summary.understandYourScore.good.text=Medelstora chanser att komma på jobbintervju
report.summary.understandYourScore.excellent.text=Mycket stor chans att komma på jobbintervju

report.analysis.title=Expert Advice


# Order Step Product Selection page

order.productSelection.title=Välj produkt
order.productSelection.subtitle=Hur kan vi hjälpa dig?
order.productSelection.submitBtn.text=Fortsätt till nästa steg
order.productSelection.validation.emptyCart=Du behöver välja minst 1 produkt för att fortsätta

order.productSelection.productsSection.title=Produkter
order.productSelection.productsSection.offerTwoProductsSameOrder.text=Spara <strong>{reductionPrice}</strong> när du beställer 2 produkter!
order.productSelection.productsSection.offerThreeProductsSameOrder.text=Spara <strong>{reductionPrice}</strong> när du beställer alla 3 produkterna!
order.productSelection.productsSection.allOffersActivated.text=Du sparar <strong>{reductionPrice}</strong>!
order.productSelection.productsSection.productName.CV_REVIEW=Granska min cv
order.productSelection.productsSection.productName.COVER_LETTER_REVIEW=Granska mitt personliga brev
order.productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Granska min LinkedIn-profil

order.productSelection.editionsSection.title=Välj version
order.productSelection.editionsSection.subtitle=Välj vilken version som passar dig bäst
order.productSelection.editionsSection.editionDescription.text.PRO=Du har några års arbetslivserfarenhet
order.productSelection.editionsSection.editionDescription.text.YOUNG_PRO=Du har jobbat mindre än 2 år, eller är student
order.productSelection.editionsSection.editionDescription.text.EXEC=Du har (eller söker) en roll med personalansvar eller verksamhetsansvar

order.productSelection.cartSection.title=Din beställning
order.productSelection.cartSection.productsHeader.products=Produkter
order.productSelection.cartSection.productsHeader.defaultPrice=Pris
order.productSelection.cartSection.coupon.label=Har du ett presentkort eller en rabattkod från någon av våra partner?
order.productSelection.cartSection.coupon.placeholder=Rabattkod
order.productSelection.cartSection.coupon.addBtn.text=Lägg till
order.productSelection.cartSection.coupon.addBtn.loadingText=Lägger till kod... 
order.productSelection.cartSection.coupon.notFoundError=Koden kunde inte hittas eller har utgått. Vänligen kontakta kundtjänst på kontakt@cruited.com
order.productSelection.cartSection.coupon.hasReachedMaxUsesError=Koden är förbrukad. Vänligen kontakta kundtjänst på kontakt@cruited.com
order.productSelection.cartSection.subTotal=Delsumma
order.productSelection.cartSection.total=Totalt att betala


# Order Step Assessment Info page *** continue translating from here

order.assessmentInfo.title=Assessment details
order.assessmentInfo.subtitle=Tell us a bit about you
order.assessmentInfo.documentsSection.title=Your documents
order.assessmentInfo.documentsSection.subtitle=This is what we will assess.
order.assessmentInfo.jobYouSearchSection.title=The job you search
order.assessmentInfo.jobYouSearchSection.subtitle=The more we know, the more we can help you. All optional information.
order.assessmentInfo.submitBtn.text=Proceed to next step
order.assessmentInfo.validation.notSignedIn=We cannot assess your LinkedIn profile unless you sign in
order.assessmentInfo.validation.jobAdUrlIncorrect=That URL looks sad :(
order.assessmentInfo.validation.customerCommentTooLong=Limited to 512 characters

order.assessmentInfo.form.browseBtn.text=Browse...
order.assessmentInfo.form.linkedinProfile.label=Your LinkedIn profile
order.assessmentInfo.form.linkedinProfile.signInBtn.text=Sign in with LinkedIn
order.assessmentInfo.form.linkedinProfile.check.step1.text=Öppna nu <a href="https://www.linkedin.com/profile/public-profile-settings?trk=prof-edit-edit-public_profile" target="blank">dina profilinställningar</a> och se till att alla kryssrutor till höger är ifyllda. De delar du inte kryssar för kommer vi inte att kunna granska.
order.assessmentInfo.form.linkedinProfile.check.step2.text=Ta en titt på <a href="https://www.linkedin.com/profile/preview?vpa=pub" target="blank">din publika profilsida</a> och se till att all information är synlig. Det du ser här är det vi kommer att bedöma.
order.assessmentInfo.form.linkedinProfile.check.checkbox.label=Klart! Min profil är redo för granskning
order.assessmentInfo.form.cvFile.label=Your CV
order.assessmentInfo.form.cvFile.placeHolder=PDF, Word, OpenOffice, RTF
order.assessmentInfo.form.coverLetterFile.label=Your cover letter
order.assessmentInfo.form.coverLetterFile.placeHolder=PDF, Word, OpenOffice, RTF
order.assessmentInfo.form.employerSought.label=Employer sought
order.assessmentInfo.form.positionSought.label=Position sought
order.assessmentInfo.form.jobAdUrl.label=URL of the job ad
order.assessmentInfo.form.customerComment.label=Do you have any specific question regarding your documents?
order.assessmentInfo.form.customerComment.description=Bör vi tänka på något särskilt i din granskning?
order.assessmentInfo.form.tos.text=I have read and accept the <a href="https://cruited.com/villkor/" target="_blank">Terms of Service</a>


# Order Step Account Creation page

order.accountCreation.title=Create your account
order.accountCreation.subtitle=Under which account do you want your assessment to be saved?
order.accountCreation.submitBtn.text=Register and continue
order.accountCreation.submitBtn.withEmailPrefix=Register with
order.accountCreation.validation.emailAlreadyRegistered=This email address is already registered. Please <a href="/login">Sign in</a>.
order.accountCreation.validation.linkedinAccountIdAlreadyRegistered=This LinkedIn account is already registered. <a href="/login">Sign in</a>.

order.accountCreation.registerWithLinkedin.switchLink.text=Prefer to register with email?
order.accountCreation.registerWithLinkedin.btn.text=Register with LinkedIn
order.accountCreation.registerWithLinkedin.email.label=Preferred email
order.accountCreation.registerWithLinkedin.validation.incorrectEmail=This email address looks incorrect

order.accountCreation.registerWithEmail.switchLink.text=Prefer to register using your LinkedIn account?
order.accountCreation.registerWithEmail.firstName.label=First name
order.accountCreation.registerWithEmail.firstName.placeholder=
order.accountCreation.registerWithEmail.emailAddress.label=Email address
order.accountCreation.registerWithEmail.emailAddress.placeholder=your@mail.com
order.accountCreation.registerWithEmail.password.label=Password
order.accountCreation.registerWithEmail.password.placeholder=5 chars minimum
order.accountCreation.registerWithEmail.validation.incorrectEmail=This email address looks incorrect
order.accountCreation.registerWithEmail.validation.passwordTooShort=Password should be at least 5 characters


# Order Step Payment page

order.payment.title=Payment
order.payment.subtitle=Please enter your card details
order.payment.submitBtn.text=Complete my order
order.payment.validation.invalidCardNumber=Invalid card number
order.payment.validation.invalidExpirationDate=Invalid expiration date
order.payment.success.text=Your payment was successful. You can access <a href="/">your dashboard</a> to see the status of your assessment.

order.payment.form.cardNumber.label=Card number
order.payment.form.cardNumber.placeholder=
order.payment.form.expires.month.label=Expires
order.payment.form.cvc.label=CVC
order.payment.form.cvc.placeholder=123
order.payment.form.cardholderName.label=Cardholder name


# Edit Order page

order.edit.saveBtn.text=Save


# Emails

email.resetPassword.subject=Nytt lösenord till Cruited
email.unpaidOrderReminder.subject=Complete your order
email.twoDaysAfterAssessmentDelivered.subject=Bara ett steg kvar till en granskning av din jobbansökan
email.orderComplete.free.subject=Granskning skapad
email.orderComplete.paid.subject=Orderbekräftelse/kvitto för beställning hos Cruited.com
email.orderComplete.paid.orderedProductsSeparator=och
