# Global

edition.name.PRO = Erfaren
edition.name.YOUNG_PRO = Ny i yrkeslivet
edition.name.EXEC = Chef
edition.name.CONSULT = Konsult
edition.name.ACADEMIA = Forskare


# Category titles

# CV
category.title.12 = Redovisa resultat och skapa trovärdighet
category.title.13 = Översiktligt och korrekt
category.title.14 = Rikta och var relevant

# Cover letter
category.title.7 = Framhäv potential
category.title.8 = Fokusera på arbetsgivaren
category.title.10 = Redovisa resultat och skapa trovärdighet
category.title.11 = Aktivt, kort och korrekt

# Linkedin profile
category.title.16 = Rikta och var relevant
category.title.17 = Skapa effekt och bygg räckvidd
category.title.18 = Översiktligt och korrekt
category.title.20 = Redovisa resultat och skapa trovärdighet


# Well Done comments

# CV
wellDone.comment.12 = Bra jobbat i denna kategori! Du har lyckats beskriva dina erfarenheter på ett bra sätt.
wellDone.comment.13 = Bra jobbat på detta område! Du har en snygg och överskådlig cv.
wellDone.comment.14 = Bra jobbat på detta område! Din cv är riktad till den tjänst du söker på ett bra sätt.

# Cover letter
wellDone.comment.7 = Bra jobbat i denna kategori! Du har lyckats framhäva din potential på ett bra sätt.
wellDone.comment.8 = Bra jobbat på detta område! Du visar att du är påläst om arbetsgivaren och varför du passar för tjänsten.
wellDone.comment.10 = Bra jobbat på detta område! Du framhäver dina egenskaper på ett bra och trovärdigt vis.
wellDone.comment.11 = Bra jobbat i denna kategori! Ditt brev är tydligt, snyggt och korrekt.

# Linkedin profile
wellDone.comment.16 = Bra jobbat på detta område! Din profil har en tydlig inriktning och du är relevant för din målgrupp.
wellDone.comment.17 = Bra jobbat på detta område! Fortsätt att bygga ditt nätverk och var aktiv på LinkedIn.
wellDone.comment.18 = Bra jobbat på detta område! Du har en tydlig och korrekt profil.
wellDone.comment.20 = Bra jobbat i denna kategori! Din profil ger ett trovärdigt intryck och du har beskrivit dina erfarenheter och utbildningar väl.


# Report preview page

report.title = Din bedömningsrapport
report.subtitle = Bedömning
report.orderCreationDate.label = Skapad
report.tabName.cv = Bedömning av CV
report.tabName.coverLetter = Bedömning av personligt brev
report.tabName.linkedinProfile = Bedömning av LinkedIn
report.tabNameSmallScreen.cv = CV
report.tabNameSmallScreen.coverLetter = Personligt brev
report.tabNameSmallScreen.linkedinProfile = LinkedIn
report.unorderedAssessment.text = Du har inte beställt den är produkten. Du behöver göra en ny beställning för att komma åt den här produkten.
report.unorderedAssessment.orderBtn.text = Beställ en ny bedömning
