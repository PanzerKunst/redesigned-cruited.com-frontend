# Global

signIn=Sign in

product.name.CV_REVIEW=CV [Resume]
product.name.COVER_LETTER_REVIEW=Cover Letter
product.name.LINKEDIN_PROFILE_REVIEW=Linkedin Profile

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive

reduction.name.2_PRODUCTS_SAME_ORDER=2-item
reduction.name.3_PRODUCTS_SAME_ORDER=3-item


# Product selection page

productSelection.title=Product Selection
productSelection.subtitle=How can we help you?
productSelection.nextStepBtn.text=Proceed to next step

productSelection.productsSection.title=Products
productSelection.productsSection.textOfferTwoProductsSameOrder=Save <strong>{reductionPrice}</strong> off your order when you select 2 items!
productSelection.productsSection.textOfferThreeProductsSameOrder=Save <strong>{reductionPrice}</strong> off your order when you select all 3 items!
productSelection.productsSection.productName.CV_REVIEW=Review my CV
productSelection.productsSection.productName.COVER_LETTER_REVIEW=Review my Cover Letter
productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Review my Linkedin Profile

productSelection.editionsSection.title=Product Edition
productSelection.editionsSection.subtitle=Please choose which edition best suits you

productSelection.cartSection.title=Your Order
productSelection.cartSection.productsHeader.products=Products
productSelection.cartSection.productsHeader.defaultPrice=Price
productSelection.cartSection.edition=Edition
productSelection.cartSection.coupon.label=Have a valid Promotion code or a Gift Card from one of our partners?
productSelection.cartSection.coupon.field.placeholder=Coupon Code
productSelection.cartSection.coupon.addButton.text=Apply coupon
productSelection.cartSection.coupon.addButton.loadingText=Applying coupon...
productSelection.cartSection.coupon.notFoundError=Coupon not found or expired
productSelection.cartSection.subTotal=Sub-total
productSelection.cartSection.total=Total You Pay
