# Global

signIn=Sign in

product.name.CV_REVIEW=CV [Resume]
product.name.COVER_LETTER_REVIEW=Cover Letter
product.name.LINKEDIN_PROFILE_REVIEW=Linkedin Profile

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive



# Product selection page

productSelection.title=Product Selection
productSelection.subtitle=How can we help you?
productSelection.productsSection.title=Products
productSelection.productsSection.textOfferTwoProductsSameOrder=Save <strong>{reductionPrice}</strong> off your order when you select 2 items!
productSelection.productsSection.textOfferThreeProductsSameOrder=Save <strong>{reductionPrice}</strong> off your order when you select all 3 items!
productSelection.productsSection.productName.CV_REVIEW=Review my CV
productSelection.productsSection.productName.COVER_LETTER_REVIEW=Review my Cover Letter
productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Review my Linkedin Profile

productSelection.editionsSection.title=Product Edition
productSelection.editionsSection.subtitle=Please choose which edition best suits you

productSelection.cartSection.title=Your Order
productSelection.cartSection.productsHeader.products=Products
productSelection.cartSection.productsHeader.defaultPrice=Price
productSelection.cartSection.edition=Edition
