# Global

defaultAssessmentTitle=Bedömning

product.name.CV_REVIEW=Granskning av CV
product.name.COVER_LETTER_REVIEW=Granskning av personligt brev
product.name.LINKEDIN_PROFILE_REVIEW=Granskning av LinkedIn

edition.name.PRO=Erfaren
edition.name.YOUNG_PRO=Ny i yrkeslivet
edition.name.EXEC=Chef

reduction.name.2_PRODUCTS_SAME_ORDER=2 dokument
reduction.name.3_PRODUCTS_SAME_ORDER=3 dokument

order.status.label=Status
order.status.notPaid.text=Betalning saknas
order.status.paid.text=Avvaktar granskning
order.status.inProgress.text=Granskning pågår
order.status.completed.text=Granskning genomförd

order.creationDate.label=Skapad

category.CV_REVIEW.12.title=Redovisa resultat och skapa trovärdighet
category.CV_REVIEW.12.shortDesc=En cv handlar i stor utsträckning om att bekräfta sin kompetens. Det är därför mycket viktigt att redovisa de resultat man uppnått.
category.CV_REVIEW.13.title=Översiktligt och korrekt
category.CV_REVIEW.13.shortDesc=Din cv ska ge arbetsgivaren en snabb översikt över dina erfarenheter och meriter. Den ska vara korrekt skriven, kort och koncis. Det finns även ett antal faktorer i språk och upplägget som påverkar hur du uppfattas som person.
category.CV_REVIEW.14.title=Rikta och var relevant
category.CV_REVIEW.14.shortDesc=I en effektiv cv är varje del relevant för det aktuella jobbet och den aktuella arbetsgivaren. Det kräver att cvn har en tydlig röd linje och att alla delar pekar i samma riktning.
category.COVER_LETTER_REVIEW.7.title=Framhäv potential
category.COVER_LETTER_REVIEW.7.shortDesc=Fokusera mer på din potential och vad du kan åstadkomma i framtiden, än på historia och vad du gjort tidigare.
category.COVER_LETTER_REVIEW.8.title=Fokusera på arbetsgivaren
category.COVER_LETTER_REVIEW.8.shortDesc=Förklara varför du valt just den här arbetsgivaren och tjänsten.
category.COVER_LETTER_REVIEW.10.title=Redovisa resultat och skapa trovärdighet
category.COVER_LETTER_REVIEW.10.shortDesc=Visa på ett trovärdigt sätt att du har kunskapen och förmågan att åstadkomma resultat för arbetsgivaren.
category.COVER_LETTER_REVIEW.11.title=Aktivt, kort och korrekt
category.COVER_LETTER_REVIEW.11.shortDesc=En dåligt skriven ansökan placerar dig som sökande ofta direkt längst ner i högen.
category.LINKEDIN_PROFILE_REVIEW.16.title=Rikta och var relevant
category.LINKEDIN_PROFILE_REVIEW.16.shortDesc=Nyckeln till framgång bland miljontals profiler på LinkedIn är att vara relevant. Du behöver visa en röd linje, få fram en bild av vart du är på väg och vad du söker. I vår granskning tittar vi på flera faktorer som rör relevans och riktning.
category.LINKEDIN_PROFILE_REVIEW.17.title=Skapa effekt och bygg räckvidd
category.LINKEDIN_PROFILE_REVIEW.17.shortDesc=Att finnas på LinkedIn är grundläggande när man söker jobb. Men för att nå framgång med LinkedIn behöver man synas och underlätta kontaktskapande. Den här kategorin handlar om hur du lyckas skapa effekt och nå ut med din profil.
category.LINKEDIN_PROFILE_REVIEW.18.title=Översiktligt och korrekt
category.LINKEDIN_PROFILE_REVIEW.18.shortDesc=Din LinkedIn-profil ska vara korrekt skriven och lätt att ta till sig. För att bli hittad av rekryterare och andra som vill nå dig, är det också viktigt att profilen är komplett och att du fyllt i rätt uppgifter på rätt plats.
category.LINKEDIN_PROFILE_REVIEW.20.title=Redovisa resultat och skapa trovärdighet
category.LINKEDIN_PROFILE_REVIEW.20.shortDesc=LinkedIn är världens största cv-bank och att berätta om sina erfarenheter och utbildningar är grundläggande. För att få kontakter och skapa möjligheter till jobb behöver du ge trovärdig bild av din bakgrund.

reportSummary.CV_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV granskningarna är <strong>{averageScore}</strong>.
reportSummary.CV_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV granskningarna är <strong>{averageScore}</strong>.
reportSummary.CV_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV granskningarna är <strong>{averageScore}</strong>.
reportSummary.CV_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV granskningarna är <strong>{averageScore}</strong>.
reportSummary.CV_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV granskningarna är <strong>{averageScore}</strong>.
reportSummary.COVER_LETTER_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av personligt brev är <strong>{averageScore}</strong>.
reportSummary.COVER_LETTER_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av personligt brev är <strong>{averageScore}</strong>.
reportSummary.COVER_LETTER_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av personligt brev är <strong>{averageScore}</strong>.
reportSummary.COVER_LETTER_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av personligt brev är <strong>{averageScore}</strong>.
reportSummary.COVER_LETTER_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av personligt brev är <strong>{averageScore}</strong>.
reportSummary.LINKEDIN_PROFILE_REVIEW.0=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
reportSummary.LINKEDIN_PROFILE_REVIEW.25=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
reportSummary.LINKEDIN_PROFILE_REVIEW.51=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
reportSummary.LINKEDIN_PROFILE_REVIEW.74=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
reportSummary.LINKEDIN_PROFILE_REVIEW.92=Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår granskning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste granskningarna av LinkedIn-profil är <strong>{averageScore}</strong>.


# Header menu

menu.signIn=Logga in
menu.signOut=Logga ut
menu.myAccount=Mitt konto


# Footer


# Sign In page

signIn.title=Logga in
signIn.methodSeparatorText=eller
signIn.validation.incorrectEmail=Den här e-postadressen ser inte korrekt ut
signIn.validation.linkedinAccountUnregistered=Vi kunde inte hitta ett konto hos oss kopplat till ditt på LinkedIn. Du kanske registrerade dig hos oss med din e-postadress?
signIn.validation.emailNotRegistered=Vi har inget konto med den här adressen
signIn.validation.emailRegisteredPasswordNull=Du har registrerat dig med ditt LinkedIn-konto.<br />Använd LinkedIn för att logga in.
signIn.validation.emailRegisteredPasswordMismatchLinkedinNotRegistered=Felaktigt lösenord. Vänligen försök igen!
signIn.validation.emailRegisteredPasswordMismatchLinkedinRegistered=Felaktigt lösenord.<br />Vi hittade en LinkedIn-profil med den här e-postadressen, så logga gärna in med LinkedIn istället.

signIn.form.linkedIn.btn.text=Logga in med LinkedIn
signIn.form.email.emailAddress.label=E-postadress
signIn.form.email.emailAddress.placeholder=din@e-post.com
signIn.form.email.password.label=Lösenord
signin.form.email.submitBtn.text=Logga in
signIn.form.forgottenPasswordLink.text=Jag behöver ett nytt lösenord


# My Account page

myAccount.title=Mitt konto
myAccount.validation.passwordTooShort=Lösenordet behöver vara minst 5 tecken
myAccount.saveSuccessful.text=Ditt konto har uppdaterats

myAccount.form.emailAddress.label=E-postadress
myAccount.form.firstName.label=Förnamn
myAccount.form.password.label=Nytt lösenord (bara om du vill byta)
myAccount.form.password.placeholder=Minst 5 tecken
myAccount.form.submitBtn.text=Spara


# Reset password pages

resetPassword.title=Återställ ditt lösenord
resetPassword.validation.incorrectEmail=Den här e-postadressen ser inte korrekt ut
resetPassword.validation.noAccountFoundForThisEmailAddress=Vi har inget konto med den här adressen
resetPassword.emailSent.text=Vi har skickat ett mejl till dig med instruktioner om hur du återställer ditt lösenord

resetPassword.form.emailAddress.label=E-postadress
resetPassword.form.emailAddress.placeholder=din@e-post.com
resetPassword.form.submitBtn.text=Jag behöver ett nytt lösenord

resetPassword.new.saveSuccessful.text=Ditt nya lösenord är sparat. Nu kan du <a href="/login">logga in</a>.
resetPassword.new.validation.passwordTooShort=Lösenordet behöver vara minst 5 tecken
resetPassword.new.form.password.label=Nytt lösenord
resetPassword.new.form.password.placeholder=Minst 5 tecken
resetPassword.new.form.submitBtn.text=Spara


# Dashboard page

dashboard.title=Mina granskningar
dashboard.subtitle=Välkommen, {firstName}!
dashboard.orderCompleted.alert.text=Din beställning har tagits emot, tack!<br />Vi kommer att meddela dig via e-post när din granskning påbörjas.
dashboard.assessmentWaiting.alert.text=Vi kommer snart att börja med din granskning.<br />Du får ett meddelande när granskningen inleds.
dashboard.assessmentInProgress.alert.text=Vi har påbörjat din granskning!<br />Du får ett meddelande när granskningen är genomförd.
dashboard.completePaymentLink.text=Betala
dashboard.newAssessmentBtn.text=Ny granskning
dashboard.viewReportBtn.text=Visa rapport
dashboard.editOrder.text=Den här granskningen har inte påbörjats och du kan fortfarande <a href="{url}">redigera din information</a> om du vill.


# Report page

report.title=Din granskningsrapport
report.unorderedAssessment.text=Du har inte beställt den är produkten. Du behöver göra en ny beställning för att komma åt den här produkten.
report.unorderedAssessment.orderBtn.text=Beställ en ny granskning
report.tabNameSmallScreen.CV_REVIEW=CV
report.tabNameSmallScreen.COVER_LETTER_REVIEW=Personligt brev
report.tabNameSmallScreen.LINKEDIN_PROFILE_REVIEW=LinkedIn

report.summary.title=Resultat av din granskning
report.summary.documentLink.text=Original
report.summary.score.label=Din C-Score
report.summary.score.bar.label.weak=Svag
report.summary.score.bar.label.good=Bra
report.summary.score.bar.label.excellent=Utmärkt
report.summary.understandYourScore.title=Förstå din C-Score
report.summary.understandYourScore.cScoreExplanation.text=C-Score mäter hur effektiv din ansökan är på en skala från 0 till 100. <a href="https://www.cruited.com/var-metod" target="_blank">Läs mer</a>
report.summary.understandYourScore.weak.text=Mycket låg chans att komma på jobbintervju
report.summary.understandYourScore.good.text=Medelstora chanser att komma på jobbintervju
report.summary.understandYourScore.excellent.text=Mycket stor chans att komma på jobbintervju

report.analysis.title=Det här behöver du förbättra
report.analysis.explanation.text=Vi har bedömt {docLabel} och identifierat vad du kan förbättra. Vi har sammanställt de åtgärder som är viktigast för att ta vidare {docLabel}. Läs igenom alla råd och börja sen förbättra {docLabel}.
report.analysis.explanation.docLabel.CV_REVIEW=din CV
report.analysis.explanation.docLabel.COVER_LETTER_REVIEW=ditt personliga brev
report.analysis.explanation.docLabel.LINKEDIN_PROFILE_REVIEW=din LinkedIn-profil


# Order Step Product Selection page

order.productSelection.title=Välj produkt
order.productSelection.subtitle=Hur kan vi hjälpa dig?
order.productSelection.submitBtn.text=Fortsätt till nästa steg
order.productSelection.validation.emptyCart=Du behöver välja minst 1 produkt för att fortsätta

order.productSelection.productsSection.title=Produkter
order.productSelection.productsSection.offerTwoProductsSameOrder.text=Spara <strong>{reductionPrice}</strong> när du beställer 2 produkter!
order.productSelection.productsSection.offerThreeProductsSameOrder.text=Spara <strong>{reductionPrice}</strong> när du beställer alla 3 produkterna!
order.productSelection.productsSection.allOffersActivated.text=Du sparar <strong>{reductionPrice}</strong>!
order.productSelection.productsSection.productName.CV_REVIEW=Granska min cv
order.productSelection.productsSection.productName.COVER_LETTER_REVIEW=Granska mitt personliga brev
order.productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Granska min LinkedIn-profil

order.productSelection.editionsSection.title=Välj version
order.productSelection.editionsSection.subtitle=Välj vilken version som passar dig bäst
order.productSelection.editionsSection.editionDescription.text.PRO=Du har några års arbetslivserfarenhet
order.productSelection.editionsSection.editionDescription.text.YOUNG_PRO=Du har jobbat mindre än 3 år, eller är student
order.productSelection.editionsSection.editionDescription.text.EXEC=Du har (eller söker) en roll med personalansvar eller verksamhetsansvar

order.productSelection.cartSection.title=Din beställning
order.productSelection.cartSection.productsHeader.products=Produkter
order.productSelection.cartSection.productsHeader.defaultPrice=Pris
order.productSelection.cartSection.coupon.label=Har du ett presentkort eller en rabattkod från någon av våra partner?
order.productSelection.cartSection.coupon.placeholder=Rabattkod
order.productSelection.cartSection.coupon.addBtn.text=Lägg till
order.productSelection.cartSection.coupon.addBtn.loadingText=Lägger till kod...
order.productSelection.cartSection.coupon.notFoundError=Koden kunde inte hittas. Vänligen kontakta kundtjänst på kontakt@cruited.com
order.productSelection.cartSection.subTotal=Delsumma
order.productSelection.cartSection.total=Att betala


# Order Step Assessment Info page

order.assessmentInfo.title=Detaljer för din granskning
order.assessmentInfo.subtitle=Information vi behöver
order.assessmentInfo.documentsSection.title=Dina dokument
order.assessmentInfo.documentsSection.subtitle=Det här är vad vi kommer att granska.
order.assessmentInfo.jobYouSearchSection.title=Jobbet du söker
order.assessmentInfo.jobYouSearchSection.subtitle=Ju mer vi vet, desto bättre kan vi hjälpa dig. Frivilliga uppgifter.
order.assessmentInfo.submitBtn.text=Gå vidare till nästa steg
order.assessmentInfo.validation.linkedin.notSignedIn=För att vi ska kunna granska din LinkedIn-profil behöver du logga in
order.assessmentInfo.validation.linkedin.publicProfileUrlMissing=Du har inte gjort din profil offentlig ännu och vi kan därför inte granska den
order.assessmentInfo.validation.linkedin.incompleteProfile.label=Din LinkedIn-profil saknar viktig information:
order.assessmentInfo.validation.linkedin.incompleteProfile.summaryMissing=Sammanfattning (summary) av din profil
order.assessmentInfo.validation.linkedin.incompleteProfile.latestProfessionalExperienceMissing=Minst en tidigare arbetslivserfarenhet med beskrivning
order.assessmentInfo.validation.linkedin.incompleteProfile.latestProfessionalExperienceSummaryMissing=En beskrivning av din senaste arbetslivserfarenhet
order.assessmentInfo.validation.jobAdUrlIncorrect=Den adressen ser inte rätt ut :(
order.assessmentInfo.validation.customerCommentTooLong=Högst 512 tecken
order.assessmentInfo.validation.requestEntityTooLarge=Filerna får inte vara större än 10MB totalt

order.assessmentInfo.form.browseBtn.text=Bläddra...
order.assessmentInfo.form.linkedinProfile.label=Din LinkedIn-profil
order.assessmentInfo.form.linkedinProfile.signInBtn.text=Logga in med LinkedIn
order.assessmentInfo.form.linkedinProfile.check.step1.text=Öppna nu <a href="https://www.linkedin.com/profile/public-profile-settings?trk=prof-edit-edit-public_profile" target="blank">dina profilinställningar</a> och se till att alla kryssrutor till höger är ifyllda. De delar du inte kryssar för kommer vi inte att kunna granska.
order.assessmentInfo.form.linkedinProfile.check.step2.text=Ta en titt på <a href="https://www.linkedin.com/profile/preview?vpa=pub" target="blank">din publika profilsida</a> och se till att all information är synlig. Det du ser här är det vi kommer att bedöma.
order.assessmentInfo.form.linkedinProfile.check.checkbox.label=Klart! Min profil är redo för granskning
order.assessmentInfo.form.linkedinProfile.check.incompleteProfile.rereadBtn.text=Läs in igen
order.assessmentInfo.form.linkedinProfile.check.incompleteProfile.checkbox.label=Jag förstår att min granskning kommer att bli begränsad eftersom min profil saknar viktiga delar. Fortsätt ändå.
order.assessmentInfo.form.cvFile.label=Ladda upp din cv
order.assessmentInfo.form.cvFile.placeHolder=PDF, Word, OpenOffice, RTF
order.assessmentInfo.form.coverLetterFile.label=Ditt personliga brev
order.assessmentInfo.form.coverLetterFile.placeHolder=PDF, Word, OpenOffice, RTF
order.assessmentInfo.form.employerSought.label=Arbetsgivare du söker dig till
order.assessmentInfo.form.positionSought.label=Tjänst du söker
order.assessmentInfo.form.jobAdUrl.label=Länk (url) till platsannons
order.assessmentInfo.form.customerComment.label=Har du några specifika frågor kring din granskning?
order.assessmentInfo.form.customerComment.description=Bör vi tänka på något särskilt i din granskning?
order.assessmentInfo.form.tos.text=Jag accepterar <a href="https://cruited.com/villkor/" target="_blank">användningsvillkoren</a>


# Order Step Account Creation page

order.accountCreation.title=Skapa ditt konto
order.accountCreation.subtitle=På vilket konto vill du spara din granskning?
order.accountCreation.submitBtn.text=Registrera och gå vidare
order.accountCreation.submitBtn.withEmailPrefix=Registrera med
order.accountCreation.validation.emailAlreadyRegistered=Det finns redan ett konto med den här adressen. <a href="/login">Logga in</a>.
order.accountCreation.validation.linkedinAccountIdAlreadyRegistered=Du är redan registrerad med LinkedIn. <a href="/login">Logga in</a>.

order.accountCreation.registerWithLinkedin.switch.question=Vill du hellre registrera
order.accountCreation.registerWithLinkedin.switch.link.text=med e-post
order.accountCreation.registerWithLinkedin.btn.text=Registrera med LinkedIn
order.accountCreation.registerWithLinkedin.profile.label=LinkedIn-profil
order.accountCreation.registerWithLinkedin.email.label=Använd den här e-postadressen
order.accountCreation.registerWithLinkedin.validation.incorrectEmail=Den här adressen ser inte korrekt ut

order.accountCreation.registerWithEmail.switch.question=Vill du hellre registrera
order.accountCreation.registerWithEmail.switch.link.text=med ditt LinkedIn-konto
order.accountCreation.registerWithEmail.firstName.label=Förnamn
order.accountCreation.registerWithEmail.firstName.placeholder=
order.accountCreation.registerWithEmail.emailAddress.label=E-postadress
order.accountCreation.registerWithEmail.emailAddress.placeholder=din@e-post.com
order.accountCreation.registerWithEmail.password.label=Lösenord
order.accountCreation.registerWithEmail.password.placeholder=Minst 5 tecken
order.accountCreation.registerWithEmail.validation.incorrectEmail=Den här e-postadressen ser inte korrekt ut
order.accountCreation.registerWithEmail.validation.passwordTooShort=Lösenordet behöver vara minst 5 tecken


# Order Step Payment page

order.payment.title=Betalning
order.payment.subtitle=Ange dina betaluppgifter
order.payment.submitBtn.text=Genomför beställning
order.payment.validation.invalidCardNumber=Ogiltigt kortnummer
order.payment.validation.invalidExpirationDate=Ogiltigt utgångsdatum

order.payment.form.cardNumber.label=Kortnummer
order.payment.form.cardNumber.placeholder=
order.payment.form.expires.month.label=Utgångsdatum
order.payment.form.cvc.label=CVC
order.payment.form.cvc.placeholder=123
order.payment.form.cardholderName.label=Kortinnehavarens namn


# Edit Order page

order.edit.saveBtn.text=Spara


# Emails

email.resetPassword.subject=Nytt lösenord till Cruited
email.unpaidOrderReminder.subject=Färdigställ din beställning
email.twoDaysAfterAssessmentDelivered.subject=Ett personligt råd om din granskning
email.orderComplete.free.subject=Granskning skapad
email.orderComplete.paid.subject=Orderbekräftelse/kvitto för beställning hos Cruited.com
email.orderComplete.paid.orderedProductsSeparator=och
