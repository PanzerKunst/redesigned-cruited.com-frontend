# Global

edition.name.PRO = Erfaren
edition.name.YOUNG_PRO = Ny i yrkeslivet
edition.name.EXEC = Chef
edition.name.CONSULT = Konsult
edition.name.ACADEMIA = Forskare


# Category titles

# CV
category.title.12 = Redovisa resultat och skapa trovärdighet
category.shortDesc.12 = En cv handlar i stor utsträckning om att bekräfta sin kompetens. Det är därför mycket viktigt att redovisa de resultat man uppnått.
category.title.13 = Översiktligt och korrekt
category.shortDesc.13 = Din cv ska ge arbetsgivaren en snabb översikt över dina erfarenheter och meriter. Den ska vara korrekt skriven, kort och koncis. Det finns även ett antal faktorer i språk och upplägget som påverkar hur du uppfattas som person.
category.title.14 = Rikta och var relevant
category.shortDesc.14 = I en effektiv cv är varje del relevant för det aktuella jobbet och den aktuella arbetsgivaren. Det kräver att cvn har en tydlig röd linje och att alla delar pekar i samma riktning.

# Cover letter
category.title.7 = Framhäv potential
category.shortDesc.7 = Fokusera mer på din potential och vad du kan åstadkomma i framtiden, än på historia och vad du gjort tidigare.
category.title.8 = Fokusera på arbetsgivaren
category.shortDesc.8 = Förklara varför du valt just den här arbetsgivaren och tjänsten.
category.title.10 = Redovisa resultat och skapa trovärdighet
category.shortDesc.10 = Visa på ett trovärdigt sätt att du har kunskapen och förmågan att åstadkomma resultat för arbetsgivaren.
category.title.11 = Aktivt, kort och korrekt
category.shortDesc.11 = En dåligt skriven ansökan placerar dig som sökande ofta direkt längst ner i högen.

# Linkedin profile
category.title.16 = Rikta och var relevant
category.shortDesc.16 = Nyckeln till framgång bland miljontals profiler på LinkedIn är att vara relevant. Du behöver visa en röd linje, få fram en bild av vart du är på väg och vad du söker. I vår bedömning tittar vi på flera faktorer som rör relevans och riktning.
category.title.17 = Skapa effekt och bygg räckvidd
category.shortDesc.17 = Att finnas på LinkedIn är grundläggande när man söker jobb. Men för att nå framgång med LinkedIn behöver man synas och underlätta kontaktskapande. Den här kategorin handlar om hur du lyckas skapa effekt och nå ut med din profil.
category.title.18 = Översiktligt och korrekt
category.shortDesc.18 = Din LinkedIn-profil ska vara korrekt skriven och lätt att ta till sig. För att bli hittad av rekryterare och andra som vill nå dig, är det också viktigt att profilen är komplett och att du fyllt i rätt uppgifter på rätt plats.
category.title.20 = Redovisa resultat och skapa trovärdighet
category.shortDesc.20 = LinkedIn är världens största cv-bank och att berätta om sina erfarenheter och utbildningar är grundläggande. För att få kontakter och skapa möjligheter till jobb behöver du ge trovärdig bild av din bakgrund.


# Well Done comments

# CV
wellDone.comment.12 = Bra jobbat i denna kategori! Du har lyckats beskriva dina erfarenheter på ett bra sätt.
wellDone.comment.13 = Bra jobbat på detta område! Du har en snygg och överskådlig cv.
wellDone.comment.14 = Bra jobbat på detta område! Din cv är riktad till den tjänst du söker på ett bra sätt.

# Cover letter
wellDone.comment.7 = Bra jobbat i denna kategori! Du har lyckats framhäva din potential på ett bra sätt.
wellDone.comment.8 = Bra jobbat på detta område! Du visar att du är påläst om arbetsgivaren och varför du passar för tjänsten.
wellDone.comment.10 = Bra jobbat på detta område! Du framhäver dina egenskaper på ett bra och trovärdigt vis.
wellDone.comment.11 = Bra jobbat i denna kategori! Ditt brev är tydligt, snyggt och korrekt.

# Linkedin profile
wellDone.comment.16 = Bra jobbat på detta område! Din profil har en tydlig inriktning och du är relevant för din målgrupp.
wellDone.comment.17 = Bra jobbat på detta område! Fortsätt att bygga ditt nätverk och var aktiv på LinkedIn.
wellDone.comment.18 = Bra jobbat på detta område! Du har en tydlig och korrekt profil.
wellDone.comment.20 = Bra jobbat i denna kategori! Din profil ger ett trovärdigt intryck och du har beskrivit dina erfarenheter och utbildningar väl.


# Report preview page

report.title = Din bedömningsrapport
report.subtitle = Bedömning
report.orderCreationDate.label = Skapad
report.tabName.cv = Bedömning av CV
report.tabName.coverLetter = Bedömning av personligt brev
report.tabName.linkedinProfile = Bedömning av LinkedIn
report.tabNameSmallScreen.cv = CV
report.tabNameSmallScreen.coverLetter = Personligt brev
report.tabNameSmallScreen.linkedinProfile = LinkedIn
report.unorderedAssessment.text = Du har inte beställt den är produkten. Du behöver göra en ny beställning för att komma åt den här produkten.
report.unorderedAssessment.orderBtn.text = Beställ en ny bedömning

report.summary.title = Resultat av din bedömning
report.summary.documentLink.text = Original
report.summary.score.label = Din C-Score
report.summary.score.bar.label.weak = Svag
report.summary.score.bar.label.good = Bra
report.summary.score.bar.label.excellent = Utmärkt
report.summary.understandYourScore.title = Förstå din C-Score
report.summary.understandYourScore.cScoreExplanation.text = C-Score mäter hur effektiv din ansökan är på en skala från 0 till 100. <a href = "https://www.cruited.com/var-metod" target = "_blank">Läs mer</a>
report.summary.understandYourScore.weak.text = Mycket låg chans att komma på jobbintervju
report.summary.understandYourScore.good.text = Medelstora chanser att komma på jobbintervju
report.summary.understandYourScore.excellent.text = Mycket stor chans att komma på jobbintervju

report.summary.cv.0 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV bedömningarna är <strong>{averageScore}</strong>.
report.summary.cv.25 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV bedömningarna är <strong>{averageScore}</strong>.
report.summary.cv.51 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV bedömningarna är <strong>{averageScore}</strong>.
report.summary.cv.74 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV bedömningarna är <strong>{averageScore}</strong>.
report.summary.cv.92 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din CV. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste CV bedömningarna är <strong>{averageScore}</strong>.
report.summary.coverLetter.0 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av personligt brev är <strong>{averageScore}</strong>.
report.summary.coverLetter.25 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av personligt brev är <strong>{averageScore}</strong>.
report.summary.coverLetter.51 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av personligt brev är <strong>{averageScore}</strong>.
report.summary.coverLetter.74 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av personligt brev är <strong>{averageScore}</strong>.
report.summary.coverLetter.92 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av ditt personliga brev. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av personligt brev är <strong>{averageScore}</strong>.
report.summary.linkedinProfile.0 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
report.summary.linkedinProfile.25 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
report.summary.linkedinProfile.51 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
report.summary.linkedinProfile.74 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av LinkedIn-profil är <strong>{averageScore}</strong>.
report.summary.linkedinProfile.92 = Du fick resultatet <strong>{score} av 100</strong> möjliga poäng i vår bedömning av din LinkedIn-profil. Genomsnittet för de {nbLastAssessmentsToTakeIntoAccount} senaste bedömningarna av LinkedIn-profil är <strong>{averageScore}</strong>.

report.analysis.title = Det här behöver du förbättra
report.analysis.explanation.text = Vi har bedömt {docLabel} och identifierat vad du kan förbättra. Vi har sammanställt de åtgärder som är viktigast för att ta vidare {docLabel}. Läs igenom alla råd och börja sen förbättra {docLabel}.
report.analysis.explanation.docLabel.cv = din CV
report.analysis.explanation.docLabel.coverLetter = ditt personliga brev
report.analysis.explanation.docLabel.linkedinProfile = din LinkedIn-profil


# Emails

email.reportAvailable.subject = Din bedömning är klar!
