# Global
signIn=Sign in

# Product selection page
productSelection.title=Product Selection
productSelection.subtitle=How can we help you?
productSelection.productsSection.title=Products
productSelection.productsSection.productName.CV_REVIEW=Review my CV
productSelection.productsSection.productName.COVER_LETTER_REVIEW=Review my Cover Letter
productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Review my Linkedin Profile
