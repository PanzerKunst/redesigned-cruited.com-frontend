home.signInWithLinkedIn=Logga in med Linkedin
