# Global

signIn=Sign in

product.name.CV_REVIEW=CV [Resume]
product.name.COVER_LETTER_REVIEW=Cover Letter
product.name.LINKEDIN_PROFILE_REVIEW=Linkedin Profile

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive

reduction.name.2_PRODUCTS_SAME_ORDER=2-item
reduction.name.3_PRODUCTS_SAME_ORDER=3-item


# Order Step Product Selection page

order.productSelection.title=Product Selection
order.productSelection.subtitle=How can we help you?
order.productSelection.nextStepBtn.text=Proceed to next step

order.productSelection.productsSection.title=Products
order.productSelection.productsSection.offerTwoProductsSameOrder.text=Save <strong>{reductionPrice}</strong> off your order when you select 2 items!
order.productSelection.productsSection.offerThreeProductsSameOrder.text=Save <strong>{reductionPrice}</strong> off your order when you select all 3 items!
order.productSelection.productsSection.productName.CV_REVIEW=Review my CV
order.productSelection.productsSection.productName.COVER_LETTER_REVIEW=Review my Cover Letter
order.productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Review my Linkedin Profile

order.productSelection.editionsSection.title=Product Edition
order.productSelection.editionsSection.subtitle=Please choose which edition best suits you

order.productSelection.cartSection.title=Your Order
order.productSelection.cartSection.productsHeader.products=Products
order.productSelection.cartSection.productsHeader.defaultPrice=Price
order.productSelection.cartSection.edition=Edition
order.productSelection.cartSection.coupon.label=Have a valid Promotion code or a Gift Card from one of our partners?
order.productSelection.cartSection.coupon.field.placeholder=Coupon Code
order.productSelection.cartSection.coupon.addBtn.text=Apply coupon
order.productSelection.cartSection.coupon.addBtn.loadingText=Applying coupon...
order.productSelection.cartSection.coupon.notFoundError=Coupon not found or expired
order.productSelection.cartSection.subTotal=Sub-total
order.productSelection.cartSection.total=Total You Pay


# Order Step Assessment Info page

order.assessmentInfo.title=Assessment details
order.assessmentInfo.subtitle=Tell us a bit about you
order.assessmentInfo.nextStepBtn.text=Proceed to next step

order.assessmentInfo.form.browseBtn.text=Browse...
order.assessmentInfo.form.linkedinProfile.label=Your Linkedin profile
order.assessmentInfo.form.linkedinProfile.signInBtn.text=Sign in with Linkedin
order.assessmentInfo.form.linkedinProfile.check.step1.text=Öppna nu <a href="https://www.linkedin.com/profile/public-profile-settings?trk=prof-edit-edit-public_profile" target="blank">dina profilinställningar</a> och se till att alla kryssrutor till höger är ifyllda. De delar du inte kryssar för kommer vi inte att kunna granska.
order.assessmentInfo.form.linkedinProfile.check.step2.text=Ta en titt på <a href="https://www.linkedin.com/profile/preview?vpa=pub" target="blank">din publika profilsida</a> och se till att all information är synlig. Det du ser här är det vi kommer att bedöma.
order.assessmentInfo.form.linkedinProfile.check.checkbox.label=Klart! Min profil är redo för granskning
order.assessmentInfo.form.linkedinProfile.validation.notSignedIn=We cannot assess your Linkedin profile unless you sign in
order.assessmentInfo.form.cvFile.label=Your CV
order.assessmentInfo.form.cvFile.placeHolder=PDF, Word, ...
order.assessmentInfo.form.coverLetterFile.label=Your cover letter
order.assessmentInfo.form.coverLetterFile.placeHolder=PDF, Word, ...
order.assessmentInfo.form.employerSought.label=Employer sought
order.assessmentInfo.form.positionSought.label=Position sought
order.assessmentInfo.form.jobAdUrl.label=URL of the job ad
order.assessmentInfo.form.tos.text=I have read and accept the <a>Terms of Service</a>


# Order Step Account Creation page

order.accountCreation.title=Create your account
order.accountCreation.subtitle=Save your order
order.accountCreation.nextStepBtn.text=Register and continue

# order.accountCreation.registerWithLinkedin.btn.text=Register with Linkedin
order.accountCreation.registerWithLinkedin.checkbox.label=Register with Linkedin
order.accountCreation.registerWithLinkedin.email.label=Preferred email
# order.accountCreation.registerWithLinkedin.validation.notSignedIn=You need to sign in if you want to register with Linkedin

order.accountCreation.registerWithEmail.checkbox.label=Register with email
order.accountCreation.registerWithEmail.firstName.label=First name
order.accountCreation.registerWithEmail.firstName.field.placeholder=
order.accountCreation.registerWithEmail.emailAddress.label=Email address
order.accountCreation.registerWithEmail.emailAddress.field.placeholder=your@mail.com
order.accountCreation.registerWithEmail.password.label=Password
order.accountCreation.registerWithEmail.password.field.placeholder=8 chars min
order.accountCreation.registerWithEmail.validation.incorrectEmail=This email address looks incorrect
order.accountCreation.registerWithEmail.validation.passwordTooShort=Password should be at least 8 characters
