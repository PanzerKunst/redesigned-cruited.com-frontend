home.signInWithLinkedIn=Logga in med Linkedin
products=Produkter
