# Global

signIn=Sign in

product.name.CV_REVIEW=CV [Resume]
product.name.COVER_LETTER_REVIEW=Cover Letter
product.name.LINKEDIN_PROFILE_REVIEW=Linkedin Profile

edition.name.PRO=Professional
edition.name.YOUNG_PRO=Young Professional
edition.name.EXEC=Executive

reduction.name.2_PRODUCTS_SAME_ORDER=2-item
reduction.name.3_PRODUCTS_SAME_ORDER=3-item


# Order Step 1 page

orderStep1.title=Product Selection
orderStep1.subtitle=How can we help you?
orderStep1.nextStepBtn.text=Proceed to next step

orderStep1.productsSection.title=Products
orderStep1.productsSection.offerTwoProductsSameOrder.text=Save <strong>{reductionPrice}</strong> off your order when you select 2 items!
orderStep1.productsSection.offerThreeProductsSameOrder.text=Save <strong>{reductionPrice}</strong> off your order when you select all 3 items!
orderStep1.productsSection.productName.CV_REVIEW=Review my CV
orderStep1.productsSection.productName.COVER_LETTER_REVIEW=Review my Cover Letter
orderStep1.productsSection.productName.LINKEDIN_PROFILE_REVIEW=Review my Linkedin Profile

orderStep1.editionsSection.title=Product Edition
orderStep1.editionsSection.subtitle=Please choose which edition best suits you

orderStep1.cartSection.title=Your Order
orderStep1.cartSection.productsHeader.products=Products
orderStep1.cartSection.productsHeader.defaultPrice=Price
orderStep1.cartSection.edition=Edition
orderStep1.cartSection.coupon.label=Have a valid Promotion code or a Gift Card from one of our partners?
orderStep1.cartSection.coupon.field.placeholder=Coupon Code
orderStep1.cartSection.coupon.addBtn.text=Apply coupon
orderStep1.cartSection.coupon.addBtn.loadingText=Applying coupon...
orderStep1.cartSection.coupon.notFoundError=Coupon not found or expired
orderStep1.cartSection.subTotal=Sub-total
orderStep1.cartSection.total=Total You Pay


# Order Step 2 page

orderStep2.title=Assessment details
orderStep2.subtitle=Tell us a bit about you
orderStep2.nextStepBtn.text=Proceed to next step

orderStep2.form.field.browseBtn.text=Browse...
orderStep2.form.field.linkedinProfile.label=Your Linkedin profile
orderStep2.form.field.linkedinProfile.signInBtn.text=Sign in with Linkedin
orderStep2.form.field.linkedinProfile.check.step1.text=Öppna nu <a href="https://www.linkedin.com/profile/public-profile-settings?trk=prof-edit-edit-public_profile" target="blank">dina profilinställningar</a> och se till att alla kryssrutor till höger är ifyllda. De delar du inte kryssar för kommer vi inte att kunna granska.
orderStep2.form.field.linkedinProfile.check.step2.text=Ta en titt på <a href="https://www.linkedin.com/profile/preview?vpa=pub" target="blank">din publika profilsida</a> och se till att all information är synlig. Det du ser här är det vi kommer att bedöma.
orderStep2.form.field.linkedinProfile.check.checkbox.label=Klart! Min profil är redo för granskning
orderStep2.form.field.linkedinProfile.validation.notSignedIn=We cannot assess your Linkedin profile unless you sign in
orderStep2.form.field.cvFile.label=Your CV
orderStep2.form.field.cvFile.placeHolder=PDF, Word, ...
orderStep2.form.field.coverLetterFile.label=Your cover letter
orderStep2.form.field.coverLetterFile.placeHolder=PDF, Word, ...
orderStep2.form.field.employerSought.label=Employer sought
orderStep2.form.field.positionSought.label=Position sought
orderStep2.form.field.jobAdUrl.label=URL of the job ad
orderStep2.form.tos.text=I have read and accept the <a>Terms of Service</a>
