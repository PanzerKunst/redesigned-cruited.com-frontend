home.title=Skriv kraftigare jobbansökningar för att få ett bättre jobb
home.subtitle=Vi granskar ditt personliga brev, CV och LinkedIn-profil. <strong>Från 299 SEK</strong>
home.hero.callToActionBtn=Kom Igång Idag
home.moneyBackGuarantee=Du omfattas av vår pengarna-tillbaka-garanti