# Global

defaultAssessmentTitle=

product.name.CV_REVIEW=
product.name.COVER_LETTER_REVIEW=
product.name.LINKEDIN_PROFILE_REVIEW=

edition.name.PRO=
edition.name.YOUNG_PRO=
edition.name.EXEC=
edition.name.short.PRO=
edition.name.short.YOUNG_PRO=
edition.name.short.EXEC=

reduction.name.2_PRODUCTS_SAME_ORDER=
reduction.name.3_PRODUCTS_SAME_ORDER=

order.status.label=
order.status.notPaid.text=
order.status.paid.text=
order.status.inProgress.text=
order.status.completed.text=

order.creationDate.label=

category.CV_REVIEW.12.title=
category.CV_REVIEW.12.shortDesc=
category.CV_REVIEW.13.title=
category.CV_REVIEW.13.shortDesc=
category.CV_REVIEW.14.title=
category.CV_REVIEW.14.shortDesc=
category.COVER_LETTER_REVIEW.7.title=
category.COVER_LETTER_REVIEW.7.shortDesc=
category.COVER_LETTER_REVIEW.8.title=
category.COVER_LETTER_REVIEW.8.shortDesc=
category.COVER_LETTER_REVIEW.10.title=
category.COVER_LETTER_REVIEW.10.shortDesc=
category.COVER_LETTER_REVIEW.11.title=
category.COVER_LETTER_REVIEW.11.shortDesc=
category.LINKEDIN_PROFILE_REVIEW.16.title=
category.LINKEDIN_PROFILE_REVIEW.16.shortDesc=
category.LINKEDIN_PROFILE_REVIEW.17.title=
category.LINKEDIN_PROFILE_REVIEW.17.shortDesc=
category.LINKEDIN_PROFILE_REVIEW.18.title=
category.LINKEDIN_PROFILE_REVIEW.18.shortDesc=
category.LINKEDIN_PROFILE_REVIEW.20.title=
category.LINKEDIN_PROFILE_REVIEW.20.shortDesc=

reportSummary.CV_REVIEW.0=
reportSummary.CV_REVIEW.25=
reportSummary.CV_REVIEW.51=
reportSummary.CV_REVIEW.74=
reportSummary.CV_REVIEW.92=
reportSummary.COVER_LETTER_REVIEW.0=
reportSummary.COVER_LETTER_REVIEW.25=
reportSummary.COVER_LETTER_REVIEW.51=
reportSummary.COVER_LETTER_REVIEW.74=
reportSummary.COVER_LETTER_REVIEW.92=
reportSummary.LINKEDIN_PROFILE_REVIEW.0=
reportSummary.LINKEDIN_PROFILE_REVIEW.25=
reportSummary.LINKEDIN_PROFILE_REVIEW.51=
reportSummary.LINKEDIN_PROFILE_REVIEW.74=
reportSummary.LINKEDIN_PROFILE_REVIEW.92=


# Header menu

menu.signIn=
menu.signOut=
menu.myAccount=


# Sign In page

signIn.title=
signIn.methodSeparatorText=
signIn.validation.incorrectEmail=
signIn.validation.invalidCredentials=
signIn.validation.linkedinAccountUnregistered=

signIn.form.linkedIn.btn.text=
signIn.form.email.emailAddress.label=
signIn.form.email.emailAddress.placeholder=
signIn.form.email.password.label=
signin.form.email.submitBtn.text=
signIn.form.forgottenPasswordLink.text=


# My Account page

myAccount.title=
myAccount.validation.passwordTooShort=
myAccount.saveSuccessful.text=

myAccount.form.emailAddress.label=
myAccount.form.firstName.label=
myAccount.form.password.label=
myAccount.form.password.placeholder=
myAccount.form.submitBtn.text=


# Reset password pages

resetPassword.title=
resetPassword.validation.incorrectEmail=
resetPassword.validation.noAccountFoundForThisEmailAddress=
resetPassword.emailSent.text=

resetPassword.form.emailAddress.label=
resetPassword.form.emailAddress.placeholder=
resetPassword.form.submitBtn.text=

resetPassword.new.saveSuccessful.text=
resetPassword.new.validation.passwordTooShort=
resetPassword.new.form.password.label=
resetPassword.new.form.password.placeholder=
resetPassword.new.form.submitBtn.text=


# Dashboard page

dashboard.title=
dashboard.subtitle=
dashboard.completePaymentLink.text=
dashboard.newAssessmentBtn.text=
dashboard.viewReportBtn.text=
dashboard.editOrder.text=


# Report page

report.title=
report.unorderedAssessment.text=
report.unorderedAssessment.orderBtn.text=

report.summary.title=
report.summary.documentLink.text=
report.summary.score.label=
report.summary.score.bar.label.weak=
report.summary.score.bar.label.good=
report.summary.score.bar.label.excellent=
report.summary.understandYourScore.title=
report.summary.understandYourScore.cScoreExplanation.text=
report.summary.understandYourScore.weak.text=
report.summary.understandYourScore.good.text=
report.summary.understandYourScore.excellent.text=

report.analysis.title=


# Order Step Product Selection page

order.productSelection.title=
order.productSelection.subtitle=
order.productSelection.submitBtn.text=
order.productSelection.validation.emptyCart=

order.productSelection.productsSection.title=
order.productSelection.productsSection.offerTwoProductsSameOrder.text=
order.productSelection.productsSection.offerThreeProductsSameOrder.text=
order.productSelection.productsSection.allOffersActivated.text=
order.productSelection.productsSection.productName.CV_REVIEW=
order.productSelection.productsSection.productName.COVER_LETTER_REVIEW=
order.productSelection.productsSection.productName.LINKEDIN_PROFILE_REVIEW=

order.productSelection.editionsSection.title=
order.productSelection.editionsSection.subtitle=
order.productSelection.editionsSection.editionDescription.text.PRO=
order.productSelection.editionsSection.editionDescription.text.YOUNG_PRO=
order.productSelection.editionsSection.editionDescription.text.EXEC=

order.productSelection.cartSection.title=
order.productSelection.cartSection.productsHeader.products=
order.productSelection.cartSection.productsHeader.defaultPrice=
order.productSelection.cartSection.coupon.label=
order.productSelection.cartSection.coupon.placeholder=
order.productSelection.cartSection.coupon.addBtn.text=
order.productSelection.cartSection.coupon.addBtn.loadingText=
order.productSelection.cartSection.coupon.notFoundError=
order.productSelection.cartSection.coupon.hasReachedMaxUsesError=
order.productSelection.cartSection.subTotal=
order.productSelection.cartSection.total=


# Order Step Assessment Info page

order.assessmentInfo.title=
order.assessmentInfo.subtitle=
order.assessmentInfo.documentsSection.title=
order.assessmentInfo.documentsSection.subtitle=
order.assessmentInfo.jobYouSearchSection.title=
order.assessmentInfo.jobYouSearchSection.subtitle=
order.assessmentInfo.submitBtn.text=
order.assessmentInfo.validation.notSignedIn=
order.assessmentInfo.validation.jobAdUrlIncorrect=
order.assessmentInfo.validation.customerCommentTooLong=

order.assessmentInfo.form.browseBtn.text=
order.assessmentInfo.form.linkedinProfile.label=
order.assessmentInfo.form.linkedinProfile.signInBtn.text=
order.assessmentInfo.form.linkedinProfile.check.step1.text=
order.assessmentInfo.form.linkedinProfile.check.step2.text=
order.assessmentInfo.form.linkedinProfile.check.checkbox.label=
order.assessmentInfo.form.cvFile.label=
order.assessmentInfo.form.cvFile.placeHolder=
order.assessmentInfo.form.coverLetterFile.label=
order.assessmentInfo.form.coverLetterFile.placeHolder=
order.assessmentInfo.form.employerSought.label=
order.assessmentInfo.form.positionSought.label=
order.assessmentInfo.form.jobAdUrl.label=
order.assessmentInfo.form.customerComment.label=
order.assessmentInfo.form.customerComment.description=
order.assessmentInfo.form.tos.text=


# Order Step Account Creation page

order.accountCreation.title=
order.accountCreation.subtitle=
order.accountCreation.submitBtn.text=
order.accountCreation.submitBtn.withEmailPrefix=
order.accountCreation.validation.emailAlreadyRegistered=
order.accountCreation.validation.linkedinAccountIdAlreadyRegistered=

order.accountCreation.registerWithLinkedin.switchLink.text=
order.accountCreation.registerWithLinkedin.btn.text=
order.accountCreation.registerWithLinkedin.email.label=
order.accountCreation.registerWithLinkedin.validation.incorrectEmail=

order.accountCreation.registerWithEmail.switchLink.text=
order.accountCreation.registerWithEmail.firstName.label=
order.accountCreation.registerWithEmail.firstName.placeholder=
order.accountCreation.registerWithEmail.emailAddress.label=
order.accountCreation.registerWithEmail.emailAddress.placeholder=
order.accountCreation.registerWithEmail.password.label=
order.accountCreation.registerWithEmail.password.placeholder=
order.accountCreation.registerWithEmail.validation.incorrectEmail=
order.accountCreation.registerWithEmail.validation.passwordTooShort=


# Order Step Payment page

order.payment.title=
order.payment.subtitle=
order.payment.submitBtn.text=
order.payment.validation.invalidCardNumber=
order.payment.validation.invalidExpirationDate=
order.payment.success.text=

order.payment.form.cardNumber.label=
order.payment.form.cardNumber.placeholder=
order.payment.form.expires.month.label=
order.payment.form.cvc.label=
order.payment.form.cvc.placeholder=
order.payment.form.cardholderName.label=


# Edit Order page

order.edit.saveBtn.text=


# Emails

email.resetPassword.subject=
email.unpaidOrderReminder.subject=
email.twoDaysAfterAssessmentDelivered.subject=
email.orderComplete.free.subject=
email.orderComplete.paid.subject=
email.orderComplete.paid.orderedProductsSeparator=